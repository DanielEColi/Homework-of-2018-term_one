----------------------------------------------------------------------------------------------------------
--ģ������: adder
--ժҪ��ʾ: 
--��ǰ�汾: 1.0.0
--ģ������: 
--�������: 20XX��XX��XX�� 
--������Ҫ:
--��Ҫע��:                                                                   
----------------------------------------------------------------------------------------------------------
--ȡ���汾: 
--ģ������:
--�������: 
--�޸�����:
--�޸��ļ�: 
----------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

---------------------------------------ENTITY DECLARATION-------------------------------------------------

entity adder is
  port(
    a_i     : in  std_logic_vector(1 downto 0);
    b_i     : in  std_logic_vector(1 downto 0);
    cin_i   : in  std_logic;
    
    sum_o   : out std_logic_vector(1 downto 0);
    cout_o  : out std_logic
    );
end adder;

----------------------------------------------------------------------------------------------------------

---------------------------------------ARCHITECTURE STRUCTURAL--------------------------------------------

architecture rtl of adder is

  signal s_carry  :  std_logic_vector(2 downto 0);
begin

  s_carry(0) <= cin_i;
  
  s_carry(1) <= (a_i(0) and b_i(0)) or (a_i(0) and s_carry(0)) or (b_i(0) and s_carry(0));
  sum_o(0) <= a_i(0) xor b_i(0) xor s_carry(0);
  
  s_carry(2) <= (a_i(1) and b_i(1)) or (a_i(1) and s_carry(1)) or (b_i(1) and s_carry(1));
  sum_o(1) <= a_i(1) xor b_i(1) xor s_carry(1);
  
  cout_o <= s_carry(2); 
end rtl;

----------------------------------------------------------------------------------------------------------
--
----------------------------------------------------------------------------------------------------------


----------------------------------------------------------------------------------------------------------
--
----------------------------------------------------------------------------------------------------------
