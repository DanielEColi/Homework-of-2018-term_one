----------------------------------------------------------------------------------------------------------
--ģ������: mux4
--ժҪ��ʾ: 
--��ǰ�汾: 1.0.0
--ģ������: 
--�������: 20XX��XX��XX�� 
--������Ҫ:
--��Ҫע��:                                                                   
----------------------------------------------------------------------------------------------------------
--ȡ���汾: 
--ģ������:
--�������: 
--�޸�����:
--�޸��ļ�: 
----------------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all; 
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

---------------------------------------ENTITY DECLARATION-------------------------------------------------
entity mux4 is
	port(
		sel : in    std_logic_vector(1 downto 0);
		y   : out 	std_logic_vector(3 downto 0)
	);
end mux4;

----------------------------------------------------------------------------------------------------------

---------------------------------------ARCHITECTURE STRUCTURAL--------------------------------------------
architecture rtl of mux4 is

begin
	process(sel)
	begin 
		case sel is
			when "00" => y <= "1110";
			when "01" => y <= "1101";
			when "10" => y <= "1011";
			when "11" => y <= "0111";
			when others => y <= "1111";
		end case;
	end process;
	
end rtl;

