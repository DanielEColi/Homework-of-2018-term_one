LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY row_scan_tb IS
END row_scan_tb;
 
ARCHITECTURE behavior OF row_scan_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT row_scan
    PORT(
         clk_i : IN  std_logic;
         rst_n_i : IN  std_logic;
         row_o : OUT  std_logic_vector(3 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal clk_i : std_logic := '0';
   signal rst_n_i : std_logic := '0';

 	--Outputs
   signal row_o : std_logic_vector(3 downto 0);

   -- Clock period definitions
   constant clk_i_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: row_scan PORT MAP (
          clk_i => clk_i,
          rst_n_i => rst_n_i,
          row_o => row_o
        );

   -- Clock process definitions
   clk_i_process :process
   begin
		clk_i <= '0';
		wait for clk_i_period/2;
		clk_i <= '1';
		wait for clk_i_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	
		rst_n_i <= '1';
      wait for clk_i_period*10;


      -- insert stimulus here 

      wait;
   end process;

END;
